module Mode_Selection(SW_SEL0, SW_SEL1, MODE);
		input SW_SEL0, SW_SEL1;
		output reg MODE;
		

endmodule
