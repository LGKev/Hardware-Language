module Top_Module_project1(SW, HEX);
	// GLOBALS
	//reg mode = 0; //maybe this is how we would select modes
	
	// INPUT

	// OUTPUT
	
	
	
	
	
	seven_segment SevenSeg0(.sw(SW), .HEX0(HEX0));
	
endmodule
